library verilog;
use verilog.vl_types.all;
entity Light_Events_vlg_vec_tst is
end Light_Events_vlg_vec_tst;
