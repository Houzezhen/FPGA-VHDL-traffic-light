library verilog;
use verilog.vl_types.all;
entity Counter_55_vlg_vec_tst is
end Counter_55_vlg_vec_tst;
