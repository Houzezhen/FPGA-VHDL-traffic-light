library verilog;
use verilog.vl_types.all;
entity Counter_0_99_vlg_vec_tst is
end Counter_0_99_vlg_vec_tst;
