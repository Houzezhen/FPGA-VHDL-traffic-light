library verilog;
use verilog.vl_types.all;
entity Block_Design_vlg_vec_tst is
end Block_Design_vlg_vec_tst;
