library verilog;
use verilog.vl_types.all;
entity Counter_5_vlg_vec_tst is
end Counter_5_vlg_vec_tst;
