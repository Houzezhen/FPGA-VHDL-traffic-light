library verilog;
use verilog.vl_types.all;
entity Road_Events_vlg_vec_tst is
end Road_Events_vlg_vec_tst;
