library verilog;
use verilog.vl_types.all;
entity COUNTER4B_vlg_vec_tst is
end COUNTER4B_vlg_vec_tst;
